module HelloWorld;
    initial
      $display ("Hello World !");
  endmodule
