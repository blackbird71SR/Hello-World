module hello_world ; #begining the module
initial begin
  $display ("Hello World by Deepak"); #print hello world
  $finish;
end
endmodule #ending the module
